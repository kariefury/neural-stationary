
*PulseLoop
.include sky130nm.lib

Xpg out2 sNoise sNoise2 sNoise sNoise sNoise sNoise sNoise2 sNoise out pg5_3
Xpg2 out sNoise sNoise2 sNoise2 sNoise2 sNoise2 sNoise2 sNoise sNoise2 out2 pg3_5


v2 sNoise  0 dc 0 trrandom (2 20p 0 0.3 0.8)
v5 sNoise2 0 dc 0 trrandom (2 20p 0 0.1 0.8)
v3 B 0 0.0
v4 VDD 0 1.8

.control
tran 1ps 35ns
plot v(out2)+4 v(out)+2 v(sNoise) v(sNoise2)-2
*hardcopy plot.ps v(out2)+4 v(out) v(sNoise)+2
*quit
.endc


*PG
.subckt pg5_3 loop A B C D E Ap Bp Cp x

xm1 1 reset_loop critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n

xm10 0 loop critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm11 Ba A critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm12 Ca B Ba 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm13 Da C Ca 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm14 Ea D Da 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm15 0 E Ea 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm16 Bpa Ap critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm17 Cpa Bp Bpa 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm18 1 Cp Cpa 1 sky130_fd_pr__pfet_01v8 l=150n w=720n

xm3 1 critical_node invO 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm4 0 critical_node invO 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm4 1 invO reset_loop 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm5 0 invO reset_loop 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm6 1 invO xe 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm7 0 invO xe 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm8 1 xe x 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm9 0 xe x 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

v1 1 0 1.8

.ends pg8

*PG
.subckt pg3_5 loop A B C Ap Bp Cp Dp Ep x

xm1 1 reset_loop critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n

xm10 0 loop critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm11 Ba A critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm12 Ca B Ba 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm13 0 C Ca 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm14 Bpa Ap critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm15 Cpa Bp Bpa 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm16 Dpa Cp Cpa 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm17 Epa Dp Dpa 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm18 1 Ep Epa 1 sky130_fd_pr__pfet_01v8 l=150n w=720n

xm3 1 critical_node invO 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm4 0 critical_node invO 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm4 1 invO reset_loop 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm5 0 invO reset_loop 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm6 1 invO xe 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm7 0 invO xe 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm8 1 xe x 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm9 0 xe x 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

v1 1 0 1.8

.ends pg3_5
