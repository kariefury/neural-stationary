magic
tech sky130A
timestamp 1632866637
<< end >>
