*PulseLoop
 .include sky130nm.lib
 Xpg sNoise out pg
 .measure tran responseTime WHEN v(out)=1.2 CROSS=1v2 sNoise 0 dc 0 trrandom (2 20p 0 0.9999999999999999 .2)
.control 
 tran 10ps 100ns 
 hardcopy plot1j v(out)+2 v(sNoise) 
quit
 .endc
 
 
 *PG
 .subckt pg A x
 
 xm1 1 reset_loop critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
 
 xm2 0 A critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
 
 xm3 1 critical_node invO 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
 xm4 0 critical_node invO 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
 
 xm4 1 invO reset_loop 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
 xm5 0 invO reset_loop 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
 
 xm6 1 invO xe 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
 xm7 0 invO xe 0 sky130_fd_pr__nfet_01v8 l=150n w=360n 
 
 xm8 1 xe x 1 sky130_fd_pr__pfet_01v8 l=150n w=720n 
 xm9 0 xe x 0 sky130_fd_pr__nfet_01v8 l=150n w=360n 
 
 
 v1 1 0 1.8 
 
 .ends pg 
 