magic
tech sky130A
timestamp 1632284168
<< nwell >>
rect -155 325 -30 420
rect -215 185 -5 325
<< nmos >>
rect -145 50 -130 150
rect -220 -125 -205 -25
<< pmos >>
rect -95 205 -80 305
<< ndiff >>
rect -195 125 -145 150
rect -195 75 -180 125
rect -160 75 -145 125
rect -195 50 -145 75
rect -130 125 -80 150
rect -130 75 -115 125
rect -95 75 -80 125
rect -130 50 -80 75
rect -270 -50 -220 -25
rect -270 -100 -255 -50
rect -235 -100 -220 -50
rect -270 -125 -220 -100
rect -205 -50 -155 -25
rect -205 -100 -190 -50
rect -170 -100 -155 -50
rect -205 -125 -155 -100
<< pdiff >>
rect -145 280 -95 305
rect -145 230 -130 280
rect -110 230 -95 280
rect -145 205 -95 230
rect -80 280 -30 305
rect -80 230 -65 280
rect -45 230 -30 280
rect -80 205 -30 230
<< ndiffc >>
rect -180 75 -160 125
rect -115 75 -95 125
rect -255 -100 -235 -50
rect -190 -100 -170 -50
<< pdiffc >>
rect -130 230 -110 280
rect -65 230 -45 280
<< psubdiff >>
rect -245 125 -195 150
rect -245 75 -225 125
rect -205 75 -195 125
rect -245 50 -195 75
rect -320 -50 -270 -25
rect -320 -100 -300 -50
rect -280 -100 -270 -50
rect -320 -125 -270 -100
<< nsubdiff >>
rect -195 280 -145 305
rect -195 230 -175 280
rect -155 230 -145 280
rect -195 205 -145 230
<< psubdiffcont >>
rect -225 75 -205 125
rect -300 -100 -280 -50
<< nsubdiffcont >>
rect -175 230 -155 280
<< poly >>
rect -120 395 -80 405
rect -120 375 -110 395
rect -90 375 -80 395
rect -120 365 -80 375
rect -95 305 -80 365
rect -95 185 -80 205
rect -145 150 -130 165
rect -145 40 -130 50
rect -145 30 -105 40
rect -145 10 -135 30
rect -115 10 -105 30
rect -145 0 -105 10
rect -220 -25 -205 -10
rect -220 -140 -205 -125
rect -220 -150 -180 -140
rect -220 -170 -210 -150
rect -190 -170 -180 -150
rect -220 -180 -180 -170
<< polycont >>
rect -110 375 -90 395
rect -135 10 -115 30
rect -210 -170 -190 -150
<< locali >>
rect -120 395 -75 405
rect -120 375 -110 395
rect -90 375 -75 395
rect -120 365 -75 375
rect -95 345 375 365
rect 355 295 375 345
rect -185 280 -105 295
rect -185 230 -175 280
rect -155 230 -130 280
rect -110 230 -105 280
rect -185 215 -105 230
rect -70 280 -40 295
rect -70 230 -65 280
rect -45 230 -40 280
rect -70 215 -40 230
rect -235 125 -155 140
rect -235 75 -225 125
rect -205 75 -180 125
rect -160 75 -155 125
rect -235 60 -155 75
rect -120 125 -90 140
rect -120 75 -115 125
rect -95 110 -90 125
rect -60 110 -40 215
rect -95 90 -40 110
rect -95 75 -90 90
rect -120 60 -90 75
rect -195 -35 -175 60
rect -145 30 -105 40
rect -145 10 -135 30
rect -115 10 -105 30
rect -60 35 -40 90
rect -60 15 -5 35
rect 10 15 20 35
rect -145 0 -105 10
rect 230 -15 250 25
rect -310 -50 -230 -35
rect -310 -100 -300 -50
rect -280 -100 -255 -50
rect -235 -100 -230 -50
rect -310 -115 -230 -100
rect -195 -50 -165 -35
rect 140 -45 160 -25
rect -195 -100 -190 -50
rect -170 -100 -165 -50
rect -195 -115 -165 -100
rect -220 -150 -180 -140
rect -220 -170 -210 -150
rect -190 -170 -180 -150
rect -220 -180 -180 -170
<< viali >>
rect -175 230 -155 280
rect -130 230 -110 280
rect -225 75 -205 125
rect -300 -100 -280 -50
rect -255 -100 -235 -50
<< metal1 >>
rect -215 280 -5 295
rect -215 230 -175 280
rect -155 230 -130 280
rect -110 230 -5 280
rect -215 220 -5 230
rect -215 215 20 220
rect 405 215 540 295
rect -310 125 105 140
rect -310 75 -225 125
rect -205 75 105 125
rect -310 60 105 75
rect -310 -50 -230 60
rect -5 45 75 60
rect -310 -100 -300 -50
rect -280 -100 -255 -50
rect -235 -100 -230 -50
rect 10 -55 75 45
rect -310 -115 -230 -100
rect -5 -70 75 -55
rect -5 -150 140 -70
rect 475 -225 540 215
rect 345 -305 540 -225
use inverter  inverter_1 /neural-stationary/Layout
timestamp 1631209646
transform 1 0 345 0 1 70
box -145 -75 60 255
use inverter  inverter_0
timestamp 1631209646
transform 1 0 140 0 1 70
box -145 -75 60 255
use inverter  inverter_2
timestamp 1631209646
transform -1 0 200 0 -1 -80
box -145 -75 60 255
use inverter  inverter_3
timestamp 1631209646
transform -1 0 -5 0 -1 -80
box -145 -75 60 255
<< labels >>
rlabel metal1 -5 255 -5 255 7 VP
rlabel locali 140 -35 140 -35 7 xe
rlabel metal1 -215 255 -215 255 7 VP
rlabel metal1 -5 100 -5 100 7 VN
rlabel space -65 -35 -65 -35 7 xout
port 3 w
rlabel metal1 489 -267 489 -267 7 Vp
port 2 w
rlabel space 142 -115 142 -115 7 VN
port 1 w
rlabel locali -135 5 -135 5 7 Ain
port 0 w
rlabel locali -220 -160 -220 -160 7 Bin
port 5 w
rlabel locali -220 -160 -220 -160 1 bin
port 6 n
<< end >>
