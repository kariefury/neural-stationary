
*PulseLoop
.include sky130nm.lib

Xpg Clk B out pg
Xpg2 out B out2 pg
Xpg3 out2 B out3 pg
Xpg4 out3 B out4 pg
Xpg5 out4 B out5 pg
Xpg6 out5 B out6 pg


*v2 Clk 0 PULSE 0 1.8 1n 20p 20p 80p 4ns
v2 Clk  0 dc 0 trrandom (2 20p 0 0.1 .8)
v3 B 0 0.0

.control
tran 0.1ns 10ns
plot v(out2)+4 v(out) v(Clk)+2
.endc


*PG
.subckt pg A B x

xm1 1 reset_loop critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n

xm2 0 A critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm10 0 B critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm3 1 critical_node invO 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm4 0 critical_node invO 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm4 1 invO reset_loop 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm5 0 invO reset_loop 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm6 1 invO xe 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm7 0 invO xe 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm8 1 xe x 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm9 0 xe x 0 sky130_fd_pr__nfet_01v8 l=150n w=360n


v1 1 0 1.8

.ends pg
