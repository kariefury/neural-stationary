
*PulseLoop
.include sky130nm.lib

Xpg out2 sNoise sNoise sNoise sNoise sNoise sNoise sNoise sNoise out pg5_3
Xpg2 out sNoise sNoise sNoise sNoise sNoise sNoise sNoise sNoise out2 pg3_5


v2 sNoise  0 dc 0 trrandom (2 20p 0 0.1 .8)
v3 B 0 0.0
v4 VDD 0 1.8

.control
tran 0.1ns 100ns
plot v(out2)+4 v(out) v(sNoise)+2
.endc


*PG
.subckt pg5_3 loop A B C D E Ap Bp Cp x

xm1 1 reset_loop critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n

xm10 0 loop critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm11 0 A critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm12 0 B critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm13 0 C critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm14 0 D critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm15 0 E critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm16 1 Ap critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm17 1 Bp critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm18 1 Cp critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm3 1 critical_node invO 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm4 0 critical_node invO 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm4 1 invO reset_loop 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm5 0 invO reset_loop 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm6 1 invO xe 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm7 0 invO xe 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm8 1 xe x 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm9 0 xe x 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

v1 1 0 1.8

.ends pg8

*PG
.subckt pg3_5 loop A B C Ap Bp Cp Dp Ep x

xm1 1 reset_loop critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n

xm10 0 loop critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm11 0 A critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm12 0 B critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm13 0 C critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm14 1 Ap critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm15 1 Bp critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm16 1 Cp critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm17 1 Dp critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm18 1 Ep critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n

xm3 1 critical_node invO 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm4 0 critical_node invO 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm4 1 invO reset_loop 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm5 0 invO reset_loop 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm6 1 invO xe 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm7 0 invO xe 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm8 1 xe x 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm9 0 xe x 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

v1 1 0 1.8

.ends pg3_5
