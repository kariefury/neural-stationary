magic
tech sky130A
timestamp 1632934578
<< nwell >>
rect -145 115 60 255
<< nmos >>
rect -25 -20 -10 80
<< pmos >>
rect -25 135 -10 235
<< ndiff >>
rect -75 55 -25 80
rect -75 5 -60 55
rect -40 5 -25 55
rect -75 -20 -25 5
rect -10 55 40 80
rect -10 5 5 55
rect 25 5 40 55
rect -10 -20 40 5
<< pdiff >>
rect -75 210 -25 235
rect -75 160 -60 210
rect -40 160 -25 210
rect -75 135 -25 160
rect -10 210 40 235
rect -10 160 5 210
rect 25 160 40 210
rect -10 135 40 160
<< ndiffc >>
rect -60 5 -40 55
rect 5 5 25 55
<< pdiffc >>
rect -60 160 -40 210
rect 5 160 25 210
<< psubdiff >>
rect -125 55 -75 80
rect -125 5 -105 55
rect -85 5 -75 55
rect -125 -20 -75 5
<< nsubdiff >>
rect -125 210 -75 235
rect -125 160 -105 210
rect -85 160 -75 210
rect -125 135 -75 160
<< psubdiffcont >>
rect -105 5 -85 55
<< nsubdiffcont >>
rect -105 160 -85 210
<< poly >>
rect -25 235 -10 250
rect -25 80 -10 135
rect -25 -35 -10 -20
rect -50 -45 -10 -35
rect -50 -65 -40 -45
rect -20 -65 -10 -45
rect -50 -75 -10 -65
<< polycont >>
rect -40 -65 -20 -45
<< locali >>
rect -115 210 -35 225
rect -115 160 -105 210
rect -85 160 -60 210
rect -40 160 -35 210
rect -115 145 -35 160
rect 0 210 30 225
rect 0 160 5 210
rect 25 160 30 210
rect 0 145 30 160
rect 10 70 30 145
rect -115 55 -35 70
rect -115 5 -105 55
rect -85 5 -60 55
rect -40 5 -35 55
rect -115 -10 -35 5
rect 0 55 30 70
rect 0 5 5 55
rect 25 5 30 55
rect 0 -10 30 5
rect -145 -45 -10 -35
rect -145 -55 -40 -45
rect -50 -65 -40 -55
rect -20 -65 -10 -45
rect 10 -55 30 -10
rect -50 -75 -10 -65
<< viali >>
rect -105 160 -85 210
rect -60 160 -40 210
rect -105 5 -85 55
rect -60 5 -40 55
<< metal1 >>
rect -145 210 60 225
rect -145 160 -105 210
rect -85 160 -60 210
rect -40 160 60 210
rect -145 145 60 160
rect -145 55 60 70
rect -145 5 -105 55
rect -85 5 -60 55
rect -40 5 60 55
rect -145 -10 60 5
<< labels >>
rlabel locali -145 -45 -145 -45 7 A
port 1 w
rlabel locali 23 -33 23 -33 1 Y
port 2 n
rlabel metal1 -141 185 -141 185 3 VP
port 3 e
rlabel metal1 -138 26 -138 26 1 VN
port 4 n
<< end >>
