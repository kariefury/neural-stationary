magic
tech sky130A
timestamp 1632936747
<< nwell >>
rect -280 325 -30 420
rect -930 185 -5 325
<< nmos >>
rect -770 30 -755 130
rect -705 30 -690 130
rect -640 30 -625 130
rect -575 30 -560 130
rect -510 30 -495 130
rect -445 30 -430 130
rect -380 30 -365 130
rect -315 30 -300 130
rect -115 5 -100 105
<< pmos >>
rect -775 205 -760 305
rect -710 205 -695 305
rect -645 205 -630 305
rect -580 205 -565 305
rect -515 205 -500 305
rect -450 205 -435 305
rect -385 205 -370 305
rect -320 205 -305 305
rect -95 205 -80 305
<< ndiff >>
rect -820 105 -770 130
rect -820 55 -805 105
rect -785 55 -770 105
rect -820 30 -770 55
rect -755 105 -705 130
rect -755 55 -740 105
rect -720 55 -705 105
rect -755 30 -705 55
rect -690 105 -640 130
rect -690 55 -675 105
rect -655 55 -640 105
rect -690 30 -640 55
rect -625 105 -575 130
rect -625 55 -610 105
rect -590 55 -575 105
rect -625 30 -575 55
rect -560 105 -510 130
rect -560 55 -545 105
rect -525 55 -510 105
rect -560 30 -510 55
rect -495 105 -445 130
rect -495 55 -480 105
rect -460 55 -445 105
rect -495 30 -445 55
rect -430 105 -380 130
rect -430 55 -415 105
rect -395 55 -380 105
rect -430 30 -380 55
rect -365 105 -315 130
rect -365 55 -350 105
rect -330 55 -315 105
rect -365 30 -315 55
rect -300 105 -250 130
rect -300 55 -285 105
rect -265 55 -250 105
rect -300 30 -250 55
rect -165 80 -115 105
rect -165 30 -150 80
rect -130 30 -115 80
rect -165 5 -115 30
rect -100 80 -50 105
rect -100 30 -85 80
rect -65 30 -50 80
rect -100 5 -50 30
<< pdiff >>
rect -825 280 -775 305
rect -825 230 -810 280
rect -790 230 -775 280
rect -825 205 -775 230
rect -760 280 -710 305
rect -760 230 -745 280
rect -725 230 -710 280
rect -760 205 -710 230
rect -695 280 -645 305
rect -695 230 -680 280
rect -660 230 -645 280
rect -695 205 -645 230
rect -630 280 -580 305
rect -630 230 -615 280
rect -595 230 -580 280
rect -630 205 -580 230
rect -565 280 -515 305
rect -565 230 -550 280
rect -530 230 -515 280
rect -565 205 -515 230
rect -500 280 -450 305
rect -500 230 -485 280
rect -465 230 -450 280
rect -500 205 -450 230
rect -435 280 -385 305
rect -435 230 -420 280
rect -400 230 -385 280
rect -435 205 -385 230
rect -370 280 -320 305
rect -370 230 -355 280
rect -335 230 -320 280
rect -370 205 -320 230
rect -305 280 -255 305
rect -305 230 -290 280
rect -270 230 -255 280
rect -305 205 -255 230
rect -140 280 -95 305
rect -140 230 -130 280
rect -110 230 -95 280
rect -140 205 -95 230
rect -80 280 -30 305
rect -80 230 -65 280
rect -45 230 -30 280
rect -80 205 -30 230
<< ndiffc >>
rect -805 55 -785 105
rect -740 55 -720 105
rect -675 55 -655 105
rect -610 55 -590 105
rect -545 55 -525 105
rect -480 55 -460 105
rect -415 55 -395 105
rect -350 55 -330 105
rect -285 55 -265 105
rect -150 30 -130 80
rect -85 30 -65 80
<< pdiffc >>
rect -810 230 -790 280
rect -745 230 -725 280
rect -680 230 -660 280
rect -615 230 -595 280
rect -550 230 -530 280
rect -485 230 -465 280
rect -420 230 -400 280
rect -355 230 -335 280
rect -290 230 -270 280
rect -130 230 -110 280
rect -65 230 -45 280
<< psubdiff >>
rect -870 105 -820 130
rect -870 55 -850 105
rect -830 55 -820 105
rect -870 30 -820 55
rect -215 80 -165 105
rect -215 30 -195 80
rect -175 30 -165 80
rect -215 5 -165 30
<< nsubdiff >>
rect -875 280 -825 305
rect -875 230 -855 280
rect -835 230 -825 280
rect -875 205 -825 230
rect -190 280 -140 305
rect -190 230 -170 280
rect -150 230 -140 280
rect -190 205 -140 230
<< psubdiffcont >>
rect -850 55 -830 105
rect -195 30 -175 80
<< nsubdiffcont >>
rect -855 230 -835 280
rect -170 230 -150 280
<< poly >>
rect -120 395 -80 405
rect -800 380 -760 390
rect -800 360 -790 380
rect -770 360 -760 380
rect -800 350 -760 360
rect -735 380 -695 390
rect -735 360 -725 380
rect -705 360 -695 380
rect -735 350 -695 360
rect -670 380 -630 390
rect -670 360 -660 380
rect -640 360 -630 380
rect -670 350 -630 360
rect -605 380 -565 390
rect -605 360 -595 380
rect -575 360 -565 380
rect -605 350 -565 360
rect -540 380 -500 390
rect -540 360 -530 380
rect -510 360 -500 380
rect -540 350 -500 360
rect -475 380 -435 390
rect -475 360 -465 380
rect -445 360 -435 380
rect -475 350 -435 360
rect -410 380 -370 390
rect -410 360 -400 380
rect -380 360 -370 380
rect -410 350 -370 360
rect -345 380 -305 390
rect -345 360 -335 380
rect -315 360 -305 380
rect -120 375 -110 395
rect -90 375 -80 395
rect -120 365 -80 375
rect -345 350 -305 360
rect -775 305 -760 350
rect -710 305 -695 350
rect -645 305 -630 350
rect -580 305 -565 350
rect -515 305 -500 350
rect -450 305 -435 350
rect -385 305 -370 350
rect -320 305 -305 350
rect -95 305 -80 365
rect -775 185 -760 205
rect -710 185 -695 205
rect -645 185 -630 205
rect -580 185 -565 205
rect -515 185 -500 205
rect -450 185 -435 205
rect -385 185 -370 205
rect -320 185 -305 205
rect -95 185 -80 205
rect -770 130 -755 145
rect -705 130 -690 145
rect -640 130 -625 145
rect -575 130 -560 145
rect -510 130 -495 145
rect -445 130 -430 145
rect -380 130 -365 145
rect -315 130 -300 145
rect -115 105 -100 120
rect -770 20 -755 30
rect -705 20 -690 30
rect -640 20 -625 30
rect -575 20 -560 30
rect -510 20 -495 30
rect -445 20 -430 30
rect -380 20 -365 30
rect -315 20 -300 30
rect -770 10 -730 20
rect -770 -10 -760 10
rect -740 -10 -730 10
rect -770 -20 -730 -10
rect -705 10 -665 20
rect -705 -10 -695 10
rect -675 -10 -665 10
rect -705 -20 -665 -10
rect -640 10 -600 20
rect -640 -10 -630 10
rect -610 -10 -600 10
rect -640 -20 -600 -10
rect -575 10 -535 20
rect -575 -10 -565 10
rect -545 -10 -535 10
rect -575 -20 -535 -10
rect -510 10 -470 20
rect -510 -10 -500 10
rect -480 -10 -470 10
rect -510 -20 -470 -10
rect -445 10 -405 20
rect -445 -10 -435 10
rect -415 -10 -405 10
rect -445 -20 -405 -10
rect -380 10 -340 20
rect -380 -10 -370 10
rect -350 -10 -340 10
rect -380 -20 -340 -10
rect -315 10 -275 20
rect -315 -10 -305 10
rect -285 -10 -275 10
rect -315 -20 -275 -10
rect -115 -20 -100 5
rect -140 -30 -100 -20
rect -140 -50 -130 -30
rect -110 -50 -100 -30
rect -140 -60 -100 -50
rect 5 -56 12 -9
<< polycont >>
rect -790 360 -770 380
rect -725 360 -705 380
rect -660 360 -640 380
rect -595 360 -575 380
rect -530 360 -510 380
rect -465 360 -445 380
rect -400 360 -380 380
rect -335 360 -315 380
rect -110 375 -90 395
rect -760 -10 -740 10
rect -695 -10 -675 10
rect -630 -10 -610 10
rect -565 -10 -545 10
rect -500 -10 -480 10
rect -435 -10 -415 10
rect -370 -10 -350 10
rect -305 -10 -285 10
rect -130 -50 -110 -30
<< locali >>
rect -120 395 -75 405
rect -800 380 -760 390
rect -800 360 -790 380
rect -770 360 -760 380
rect -800 350 -760 360
rect -735 380 -695 390
rect -735 360 -725 380
rect -705 360 -695 380
rect -735 350 -695 360
rect -670 380 -630 390
rect -670 360 -660 380
rect -640 360 -630 380
rect -670 350 -630 360
rect -605 380 -565 390
rect -605 360 -595 380
rect -575 360 -565 380
rect -605 350 -565 360
rect -540 380 -500 390
rect -540 360 -530 380
rect -510 360 -500 380
rect -540 350 -500 360
rect -475 380 -435 390
rect -475 360 -465 380
rect -445 360 -435 380
rect -475 350 -435 360
rect -410 380 -370 390
rect -410 360 -400 380
rect -380 360 -370 380
rect -410 350 -370 360
rect -345 380 -305 390
rect -345 360 -335 380
rect -315 360 -305 380
rect -120 375 -110 395
rect -90 375 -75 395
rect -120 365 -75 375
rect -345 350 -305 360
rect -95 345 375 365
rect 355 295 375 345
rect -865 280 -785 295
rect -865 230 -855 280
rect -835 230 -810 280
rect -790 230 -785 280
rect -865 215 -785 230
rect -750 280 -720 295
rect -750 230 -745 280
rect -725 230 -720 280
rect -750 215 -720 230
rect -685 280 -655 295
rect -685 230 -680 280
rect -660 230 -655 280
rect -685 215 -655 230
rect -620 280 -590 295
rect -620 230 -615 280
rect -595 230 -590 280
rect -620 215 -590 230
rect -555 280 -525 295
rect -555 230 -550 280
rect -530 230 -525 280
rect -555 215 -525 230
rect -490 280 -460 295
rect -490 230 -485 280
rect -465 230 -460 280
rect -490 215 -460 230
rect -425 280 -395 295
rect -425 230 -420 280
rect -400 230 -395 280
rect -425 215 -395 230
rect -360 280 -330 295
rect -360 230 -355 280
rect -335 230 -330 280
rect -360 215 -330 230
rect -295 280 -265 295
rect -295 230 -290 280
rect -270 230 -265 280
rect -295 215 -265 230
rect -180 280 -105 295
rect -180 230 -170 280
rect -150 230 -130 280
rect -110 230 -105 280
rect -180 215 -105 230
rect -70 280 -40 295
rect -70 230 -65 280
rect -45 230 -40 280
rect -70 215 -40 230
rect -740 185 -720 215
rect -675 185 -655 215
rect -610 185 -590 215
rect -545 185 -525 215
rect -480 185 -460 215
rect -415 185 -395 215
rect -350 185 -330 215
rect -285 185 -265 215
rect -60 185 -40 215
rect -740 165 -40 185
rect -280 140 -260 165
rect -860 105 -780 120
rect -860 55 -850 105
rect -830 55 -805 105
rect -785 55 -780 105
rect -860 40 -780 55
rect -745 105 -715 120
rect -745 55 -740 105
rect -720 55 -715 105
rect -745 40 -715 55
rect -680 105 -650 120
rect -680 55 -675 105
rect -655 55 -650 105
rect -680 40 -650 55
rect -615 105 -585 120
rect -615 55 -610 105
rect -590 55 -585 105
rect -615 40 -585 55
rect -550 105 -520 120
rect -550 55 -545 105
rect -525 55 -520 105
rect -550 40 -520 55
rect -485 105 -455 120
rect -485 55 -480 105
rect -460 55 -455 105
rect -485 40 -455 55
rect -420 105 -390 120
rect -420 55 -415 105
rect -395 55 -390 105
rect -420 40 -390 55
rect -355 105 -325 120
rect -355 55 -350 105
rect -330 55 -325 105
rect -355 40 -325 55
rect -290 105 -260 140
rect -290 55 -285 105
rect -265 55 -260 105
rect -60 95 -40 165
rect -290 40 -260 55
rect -205 80 -125 95
rect -205 30 -195 80
rect -175 30 -150 80
rect -130 30 -125 80
rect -770 10 -730 20
rect -770 -10 -760 10
rect -740 -10 -730 10
rect -770 -20 -730 -10
rect -705 10 -665 20
rect -705 -10 -695 10
rect -675 -10 -665 10
rect -705 -20 -665 -10
rect -640 10 -600 20
rect -640 -10 -630 10
rect -610 -10 -600 10
rect -640 -20 -600 -10
rect -575 10 -535 20
rect -575 -10 -565 10
rect -545 -10 -535 10
rect -575 -20 -535 -10
rect -510 10 -470 20
rect -510 -10 -500 10
rect -480 -10 -470 10
rect -510 -20 -470 -10
rect -445 10 -405 20
rect -445 -10 -435 10
rect -415 -10 -405 10
rect -445 -20 -405 -10
rect -380 10 -340 20
rect -380 -10 -370 10
rect -350 -10 -340 10
rect -380 -20 -340 -10
rect -315 10 -275 20
rect -205 15 -125 30
rect -90 80 -40 95
rect -90 30 -85 80
rect -65 35 -40 80
rect -65 30 -5 35
rect -90 15 -5 30
rect 10 15 20 35
rect 150 15 202 35
rect -315 -10 -305 10
rect -285 -10 -275 10
rect -315 -20 -275 -10
rect 230 -15 250 25
rect -140 -30 -100 -20
rect -140 -50 -130 -30
rect -110 -50 -100 -30
rect 140 -45 170 -25
rect -140 -60 -100 -50
rect -33 -195 -19 -168
<< viali >>
rect -855 230 -835 280
rect -810 230 -790 280
rect -170 230 -150 280
rect -130 230 -110 280
rect -850 55 -830 105
rect -805 55 -785 105
rect -195 30 -175 80
rect -150 30 -130 80
<< metal1 >>
rect -930 280 -5 295
rect -930 230 -855 280
rect -835 230 -810 280
rect -790 230 -170 280
rect -150 230 -130 280
rect -110 230 -5 280
rect -930 220 -5 230
rect -930 215 20 220
rect -930 105 105 140
rect -930 60 -850 105
rect -860 55 -850 60
rect -830 55 -805 105
rect -785 80 105 105
rect -785 60 -195 80
rect -785 55 -250 60
rect -860 40 -250 55
rect -215 35 -195 60
rect -205 30 -195 35
rect -175 30 -150 80
rect -130 60 105 80
rect -130 30 -50 60
rect -5 45 75 60
rect -205 15 -50 30
rect 10 -55 75 45
rect -5 -70 75 -55
rect -930 -150 -65 -70
rect -5 -150 140 -70
rect 210 -150 405 -70
rect -930 -305 -65 -225
rect 345 -305 405 -225
use inverter  inverter_1
timestamp 1632934578
transform 1 0 345 0 1 70
box -145 -75 60 255
use inverter  inverter_0
timestamp 1632934578
transform 1 0 140 0 1 70
box -145 -75 60 255
use inverter  inverter_2
timestamp 1632934578
transform -1 0 200 0 -1 -80
box -145 -75 60 255
use inverter  inverter_3
timestamp 1632934578
transform -1 0 -5 0 -1 -80
box -145 -75 60 255
<< labels >>
rlabel locali 140 -35 140 -35 7 xe
rlabel space 142 -115 142 -115 7 VN
port 3 w
rlabel metal1 -15 85 10 110 7 VN
port 15 w
rlabel locali -345 350 -305 390 7 Iin
port 14 w
rlabel locali -410 370 -410 370 7 Jin
port 16 w
rlabel locali -475 370 -475 370 7 Kin
port 17 w
rlabel locali -540 370 -540 370 7 Lin
port 18 w
rlabel locali -605 370 -605 370 1 Min
port 19 n
rlabel locali -670 370 -670 370 1 Nin
port 20 n
rlabel locali -735 370 -735 370 1 Oin
port 21 n
rlabel locali -800 370 -800 370 7 Pin
port 22 w
rlabel metal1 375 -265 375 -265 7 VP
rlabel locali -25 -180 -25 -180 7 xout
rlabel locali -305 -15 -305 -15 7 Ain
port 0 w
rlabel locali -380 0 -380 0 1 bin
port 1 n
rlabel locali -380 0 -380 0 7 Bin
port 2 w
rlabel locali -510 -20 -470 20 7 Din
port 7 w
rlabel poly -640 -20 -600 20 7 Fin
port 9 w
rlabel locali -705 -20 -665 20 3 Gin
port 10 e
rlabel locali -770 -20 -730 20 7 Hin
port 11 w
rlabel locali -445 -20 -405 20 7 Cin
port 13 w
rlabel locali -575 -20 -535 20 7 Ein
port 8 w
rlabel metal1 -260 95 -260 95 3 VN
rlabel metal1 -930 95 -930 95 3 VN
rlabel metal1 -925 255 -925 255 7 VP
port 5 w
rlabel locali 35 355 35 355 7 reset_loop
rlabel space 215 -45 215 -45 1 inv2input
rlabel locali -30 -185 -20 -175 7 xout
port 4 w
rlabel locali 175 25 175 25 1 pgnode
rlabel polycont -125 -40 -125 -40 1 n_para
port 23 n
<< end >>
