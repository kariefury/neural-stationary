// Verilog test bench for example_3_1
`timescale 1ns/100ps
`include "fiveclocks.v"

module five_clocks_tb;

  reg clk;
  wire to_clock;
  reg reset;
  reg b;
  wire m;
  wire t, tt, ttt, tttt, ttttt;
  // Instantiate design under test
  fiveclocks FC(.clk(clk),.b( b ),.reset(reset),.t(t),.tt(tt),.ttt(ttt),.tttt(tttt),.ttttt(ttttt),.m(m));

   initial begin
      $dumpfile("fiveclocks.vcd");
      $dumpvars(0, five_clocks_tb);
      b = 0;
      clk = 0;
      reset = 1; 
      display;
      clk = 1;
      
      display;
      clk = 0;
      display;
      clk = 1;
      display;
      reset = 0;
       display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  1 ; display;    
clk =  0 ; display;    
clk =  1 ; display; 
   end

  task display;
    #1 $display("clk:%0h, t:%0h, tt:%0h, ttt:%0h, tttt:%0h, ttttt:%0h, m:%0h",
      clk,t, tt, ttt,tttt,ttttt,m);
  endtask

endmodule




