magic
tech sky130A
timestamp 1632866761
<< nwell >>
rect -280 325 -30 420
rect -895 185 -5 325
<< nmos >>
rect -600 30 -585 130
rect -535 30 -520 130
rect -470 30 -455 130
rect -405 30 -390 130
rect -340 30 -325 130
rect -275 30 -260 130
rect -210 30 -195 130
rect -145 30 -130 130
<< pmos >>
rect -775 205 -760 305
rect -710 205 -695 305
rect -645 205 -630 305
rect -580 205 -565 305
rect -515 205 -500 305
rect -450 205 -435 305
rect -385 205 -370 305
rect -320 205 -305 305
rect -95 205 -80 305
<< ndiff >>
rect -650 105 -600 130
rect -650 55 -635 105
rect -615 55 -600 105
rect -650 30 -600 55
rect -585 105 -535 130
rect -585 55 -570 105
rect -550 55 -535 105
rect -585 30 -535 55
rect -520 105 -470 130
rect -520 55 -505 105
rect -485 55 -470 105
rect -520 30 -470 55
rect -455 105 -405 130
rect -455 55 -440 105
rect -420 55 -405 105
rect -455 30 -405 55
rect -390 105 -340 130
rect -390 55 -375 105
rect -355 55 -340 105
rect -390 30 -340 55
rect -325 105 -275 130
rect -325 55 -310 105
rect -290 55 -275 105
rect -325 30 -275 55
rect -260 105 -210 130
rect -260 55 -245 105
rect -225 55 -210 105
rect -260 30 -210 55
rect -195 105 -145 130
rect -195 55 -180 105
rect -160 55 -145 105
rect -195 30 -145 55
rect -130 105 -80 130
rect -130 55 -115 105
rect -95 55 -80 105
rect -130 30 -80 55
<< pdiff >>
rect -825 280 -775 305
rect -825 230 -810 280
rect -790 230 -775 280
rect -825 205 -775 230
rect -760 280 -710 305
rect -760 230 -745 280
rect -725 230 -710 280
rect -760 205 -710 230
rect -695 280 -645 305
rect -695 230 -680 280
rect -660 230 -645 280
rect -695 205 -645 230
rect -630 280 -580 305
rect -630 230 -615 280
rect -595 230 -580 280
rect -630 205 -580 230
rect -565 280 -515 305
rect -565 230 -550 280
rect -530 230 -515 280
rect -565 205 -515 230
rect -500 280 -450 305
rect -500 230 -485 280
rect -465 230 -450 280
rect -500 205 -450 230
rect -435 280 -385 305
rect -435 230 -420 280
rect -400 230 -385 280
rect -435 205 -385 230
rect -370 280 -320 305
rect -370 230 -355 280
rect -335 230 -320 280
rect -370 205 -320 230
rect -305 280 -255 305
rect -305 230 -290 280
rect -270 230 -255 280
rect -305 205 -255 230
rect -140 280 -95 305
rect -140 230 -130 280
rect -110 230 -95 280
rect -140 205 -95 230
rect -80 280 -30 305
rect -80 230 -65 280
rect -45 230 -30 280
rect -80 205 -30 230
<< ndiffc >>
rect -635 55 -615 105
rect -570 55 -550 105
rect -505 55 -485 105
rect -440 55 -420 105
rect -375 55 -355 105
rect -310 55 -290 105
rect -245 55 -225 105
rect -180 55 -160 105
rect -115 55 -95 105
<< pdiffc >>
rect -810 230 -790 280
rect -745 230 -725 280
rect -680 230 -660 280
rect -615 230 -595 280
rect -550 230 -530 280
rect -485 230 -465 280
rect -420 230 -400 280
rect -355 230 -335 280
rect -290 230 -270 280
rect -130 230 -110 280
rect -65 230 -45 280
<< psubdiff >>
rect -700 105 -650 130
rect -700 55 -680 105
rect -660 55 -650 105
rect -700 30 -650 55
<< nsubdiff >>
rect -875 280 -825 305
rect -875 230 -855 280
rect -835 230 -825 280
rect -875 205 -825 230
rect -190 280 -140 305
rect -190 230 -170 280
rect -150 230 -140 280
rect -190 205 -140 230
<< psubdiffcont >>
rect -680 55 -660 105
<< nsubdiffcont >>
rect -855 230 -835 280
rect -170 230 -150 280
<< poly >>
rect -120 395 -80 405
rect -800 380 -760 390
rect -800 360 -790 380
rect -770 360 -760 380
rect -800 350 -760 360
rect -735 380 -695 390
rect -735 360 -725 380
rect -705 360 -695 380
rect -735 350 -695 360
rect -670 380 -630 390
rect -670 360 -660 380
rect -640 360 -630 380
rect -670 350 -630 360
rect -605 380 -565 390
rect -605 360 -595 380
rect -575 360 -565 380
rect -605 350 -565 360
rect -540 380 -500 390
rect -540 360 -530 380
rect -510 360 -500 380
rect -540 350 -500 360
rect -475 380 -435 390
rect -475 360 -465 380
rect -445 360 -435 380
rect -475 350 -435 360
rect -410 380 -370 390
rect -410 360 -400 380
rect -380 360 -370 380
rect -410 350 -370 360
rect -345 380 -305 390
rect -345 360 -335 380
rect -315 360 -305 380
rect -120 375 -110 395
rect -90 375 -80 395
rect -120 365 -80 375
rect -345 350 -305 360
rect -775 305 -760 350
rect -710 305 -695 350
rect -645 305 -630 350
rect -580 305 -565 350
rect -515 305 -500 350
rect -450 305 -435 350
rect -385 305 -370 350
rect -320 305 -305 350
rect -95 305 -80 365
rect -775 185 -760 205
rect -710 185 -695 205
rect -645 185 -630 205
rect -580 185 -565 205
rect -515 185 -500 205
rect -450 185 -435 205
rect -385 185 -370 205
rect -320 185 -305 205
rect -95 185 -80 205
rect -600 130 -585 145
rect -535 130 -520 145
rect -470 130 -455 145
rect -405 130 -390 145
rect -340 130 -325 145
rect -275 130 -260 145
rect -210 130 -195 145
rect -145 130 -130 145
rect -600 20 -585 30
rect -535 20 -520 30
rect -470 20 -455 30
rect -405 20 -390 30
rect -340 20 -325 30
rect -275 20 -260 30
rect -210 20 -195 30
rect -145 20 -130 30
rect -600 10 -560 20
rect -600 -10 -590 10
rect -570 -10 -560 10
rect -600 -20 -560 -10
rect -535 10 -495 20
rect -535 -10 -525 10
rect -505 -10 -495 10
rect -535 -20 -495 -10
rect -470 10 -430 20
rect -470 -10 -460 10
rect -440 -10 -430 10
rect -470 -20 -430 -10
rect -405 10 -365 20
rect -405 -10 -395 10
rect -375 -10 -365 10
rect -405 -20 -365 -10
rect -340 10 -300 20
rect -340 -10 -330 10
rect -310 -10 -300 10
rect -340 -20 -300 -10
rect -275 10 -235 20
rect -275 -10 -265 10
rect -245 -10 -235 10
rect -275 -20 -235 -10
rect -210 10 -170 20
rect -210 -10 -200 10
rect -180 -10 -170 10
rect -210 -20 -170 -10
rect -145 10 -105 20
rect -145 -10 -135 10
rect -115 -10 -105 10
rect -145 -20 -105 -10
<< polycont >>
rect -790 360 -770 380
rect -725 360 -705 380
rect -660 360 -640 380
rect -595 360 -575 380
rect -530 360 -510 380
rect -465 360 -445 380
rect -400 360 -380 380
rect -335 360 -315 380
rect -110 375 -90 395
rect -590 -10 -570 10
rect -525 -10 -505 10
rect -460 -10 -440 10
rect -395 -10 -375 10
rect -330 -10 -310 10
rect -265 -10 -245 10
rect -200 -10 -180 10
rect -135 -10 -115 10
<< locali >>
rect -120 395 -75 405
rect -800 380 -760 390
rect -800 360 -790 380
rect -770 360 -760 380
rect -800 350 -760 360
rect -735 380 -695 390
rect -735 360 -725 380
rect -705 360 -695 380
rect -735 350 -695 360
rect -670 380 -630 390
rect -670 360 -660 380
rect -640 360 -630 380
rect -670 350 -630 360
rect -605 380 -565 390
rect -605 360 -595 380
rect -575 360 -565 380
rect -605 350 -565 360
rect -540 380 -500 390
rect -540 360 -530 380
rect -510 360 -500 380
rect -540 350 -500 360
rect -475 380 -435 390
rect -475 360 -465 380
rect -445 360 -435 380
rect -475 350 -435 360
rect -410 380 -370 390
rect -410 360 -400 380
rect -380 360 -370 380
rect -410 350 -370 360
rect -345 380 -305 390
rect -345 360 -335 380
rect -315 360 -305 380
rect -120 375 -110 395
rect -90 375 -75 395
rect -120 365 -75 375
rect -345 350 -305 360
rect -95 345 375 365
rect 355 295 375 345
rect -865 280 -785 295
rect -865 230 -855 280
rect -835 230 -810 280
rect -790 230 -785 280
rect -865 215 -785 230
rect -750 280 -720 295
rect -750 230 -745 280
rect -725 230 -720 280
rect -750 215 -720 230
rect -685 280 -655 295
rect -685 230 -680 280
rect -660 230 -655 280
rect -685 215 -655 230
rect -620 280 -590 295
rect -620 230 -615 280
rect -595 230 -590 280
rect -620 215 -590 230
rect -555 280 -525 295
rect -555 230 -550 280
rect -530 230 -525 280
rect -555 215 -525 230
rect -490 280 -460 295
rect -490 230 -485 280
rect -465 230 -460 280
rect -490 215 -460 230
rect -425 280 -395 295
rect -425 230 -420 280
rect -400 230 -395 280
rect -425 215 -395 230
rect -360 280 -330 295
rect -360 230 -355 280
rect -335 230 -330 280
rect -360 215 -330 230
rect -295 280 -265 295
rect -295 230 -290 280
rect -270 230 -265 280
rect -295 215 -265 230
rect -180 280 -105 295
rect -180 230 -170 280
rect -150 230 -130 280
rect -110 230 -105 280
rect -180 215 -105 230
rect -70 280 -40 295
rect -70 230 -65 280
rect -45 230 -40 280
rect -70 215 -40 230
rect -740 185 -720 215
rect -675 185 -655 215
rect -610 185 -590 215
rect -545 185 -525 215
rect -480 185 -460 215
rect -415 185 -395 215
rect -350 185 -330 215
rect -285 185 -265 215
rect -60 185 -40 215
rect -740 165 -40 185
rect -690 105 -610 120
rect -690 55 -680 105
rect -660 55 -635 105
rect -615 55 -610 105
rect -690 40 -610 55
rect -575 105 -545 120
rect -575 55 -570 105
rect -550 55 -545 105
rect -575 40 -545 55
rect -510 105 -480 120
rect -510 55 -505 105
rect -485 55 -480 105
rect -510 40 -480 55
rect -445 105 -415 120
rect -445 55 -440 105
rect -420 55 -415 105
rect -445 40 -415 55
rect -380 105 -350 120
rect -380 55 -375 105
rect -355 55 -350 105
rect -380 40 -350 55
rect -315 105 -285 120
rect -315 55 -310 105
rect -290 55 -285 105
rect -315 40 -285 55
rect -250 105 -220 120
rect -250 55 -245 105
rect -225 55 -220 105
rect -250 40 -220 55
rect -185 105 -155 120
rect -185 55 -180 105
rect -160 55 -155 105
rect -185 40 -155 55
rect -120 110 -90 120
rect -60 110 -40 165
rect -120 105 -40 110
rect -120 55 -115 105
rect -95 90 -40 105
rect -95 55 -90 90
rect -120 40 -90 55
rect -60 35 -40 90
rect -600 10 -560 20
rect -600 -10 -590 10
rect -570 -10 -560 10
rect -600 -20 -560 -10
rect -535 10 -495 20
rect -535 -10 -525 10
rect -505 -10 -495 10
rect -535 -20 -495 -10
rect -470 10 -430 20
rect -470 -10 -460 10
rect -440 -10 -430 10
rect -470 -20 -430 -10
rect -405 10 -365 20
rect -405 -10 -395 10
rect -375 -10 -365 10
rect -405 -20 -365 -10
rect -340 10 -300 20
rect -340 -10 -330 10
rect -310 -10 -300 10
rect -340 -20 -300 -10
rect -275 10 -235 20
rect -275 -10 -265 10
rect -245 -10 -235 10
rect -275 -20 -235 -10
rect -210 10 -170 20
rect -210 -10 -200 10
rect -180 -10 -170 10
rect -210 -20 -170 -10
rect -145 10 -105 20
rect -60 15 -5 35
rect 10 15 20 35
rect 170 15 200 35
rect -145 -10 -135 10
rect -115 -10 -105 10
rect -145 -20 -105 -10
rect 230 -15 250 25
rect 140 -45 170 -25
<< viali >>
rect -855 230 -835 280
rect -810 230 -790 280
rect -170 230 -150 280
rect -130 230 -110 280
rect -680 55 -660 105
rect -635 55 -615 105
<< metal1 >>
rect -895 280 -5 295
rect -895 230 -855 280
rect -835 230 -810 280
rect -790 230 -170 280
rect -150 230 -130 280
rect -110 230 -5 280
rect -895 220 -5 230
rect -895 215 20 220
rect -895 105 105 140
rect -895 60 -680 105
rect -690 55 -680 60
rect -660 55 -635 105
rect -615 60 105 105
rect -615 55 -80 60
rect -690 40 -80 55
rect -5 45 75 60
rect 10 -55 75 45
rect -5 -70 75 -55
rect -895 -150 -65 -70
rect -5 -150 140 -70
rect 210 -150 405 -70
rect -895 -305 -65 -225
rect 345 -305 405 -225
use inverter  inverter_3
timestamp 1632865684
transform -1 0 -5 0 -1 -80
box -145 -75 60 255
use inverter  inverter_2
timestamp 1632865684
transform -1 0 200 0 -1 -80
box -145 -75 60 255
use inverter  inverter_0
timestamp 1632865684
transform 1 0 140 0 1 70
box -145 -75 60 255
use inverter  inverter_1
timestamp 1632865684
transform 1 0 345 0 1 70
box -145 -75 60 255
<< labels >>
rlabel locali 140 -35 140 -35 7 xe
rlabel space 142 -115 142 -115 7 VN
port 3 w
rlabel locali -135 -15 -135 -15 7 Ain
port 0 w
rlabel locali -210 0 -210 0 1 bin
port 1 n
rlabel locali -210 0 -210 0 7 Bin
port 2 w
rlabel locali -340 -20 -300 20 7 Din
port 7 w
rlabel poly -470 -20 -430 20 7 Fin
port 9 w
rlabel locali -535 -20 -495 20 3 Gin
port 10 e
rlabel locali -600 -20 -560 20 7 Hin
port 11 w
rlabel locali -275 -20 -235 20 7 Cin
port 13 w
rlabel locali -405 -20 -365 20 7 Ein
port 8 w
rlabel locali -10 355 -10 355 7 reset_loop
rlabel metal1 -15 85 10 110 7 VN
port 15 w
rlabel locali -345 350 -305 390 7 Iin
port 14 w
rlabel metal1 -895 255 -895 255 7 VP
port 5 w
rlabel locali -410 370 -410 370 7 Jin
port 16 w
rlabel locali -475 370 -475 370 7 Kin
port 17 w
rlabel locali -540 370 -540 370 7 Lin
port 18 w
rlabel locali -605 370 -605 370 1 Min
port 19 n
rlabel locali -670 370 -670 370 1 Nin
port 20 n
rlabel locali -735 370 -735 370 1 Oin
port 21 n
rlabel locali -800 370 -800 370 7 Pin
port 22 w
rlabel metal1 375 -265 375 -265 7 VP
rlabel metal1 -895 95 -895 95 3 VN
rlabel space -25 -180 -25 -180 7 xout
rlabel space -35 -40 -25 -30 7 xout
port 4 w
<< end >>
