* SPICE3 file created from neuron.ext - technology: sky130A

.option scale=10000u

.subckt inverter A w_n145_115# a_n10_n20# a_n125_n20#
X0 a_n10_n20# A w_n145_115# w_n145_115# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X1 a_n10_n20# A a_n125_n20# a_n125_n20# sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
C0 w_n145_115# a_n10_n20# 0.22fF
C1 A a_n125_n20# 0.53fF
C2 a_n10_n20# a_n125_n20# 0.34fF
C3 w_n145_115# a_n125_n20# 0.59fF
.ends

.subckt pg17Input8p8n_para_1n Ain bin VP Din Ein Fin Gin Hin Cin Iin VN Jin Kin Lin
+ Min Nin Oin Pin inverter_3/a_n10_n20# xe a_n140_n60# reset_loop inverter_2/A
Xinverter_0 inverter_0/A VP inverter_2/A VN inverter
Xinverter_1 inverter_2/A VP reset_loop VN inverter
Xinverter_2 inverter_2/A VP xe VN inverter
Xinverter_3 xe VP inverter_3/a_n10_n20# VN inverter
X0 a_n560_30# Ein a_n625_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X1 inverter_0/A reset_loop VP VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X2 inverter_0/A Min inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X3 a_n755_30# Hin VN VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X4 inverter_0/A Kin inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X5 a_n690_30# Gin a_n755_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X6 inverter_0/A Iin inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X7 inverter_0/A Oin inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X8 a_n365_30# bin a_n430_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X9 inverter_0/A Ain a_n365_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X10 inverter_0/A Jin inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X11 a_n495_30# Din a_n560_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X12 inverter_0/A Pin VP VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X13 inverter_0/A Nin inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X14 a_n430_30# Cin a_n495_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X15 inverter_0/A Lin inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X16 a_n625_30# Fin a_n690_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X17 inverter_0/A a_n140_n60# VN VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
C0 Iin Jin 0.12fF
C1 Cin bin 0.10fF
C2 Gin Hin 0.10fF
C3 Din Ein 0.10fF
C4 Nin Min 0.12fF
C5 Jin Kin 0.12fF
C6 Lin Kin 0.12fF
C7 Gin Fin 0.10fF
C8 VP reset_loop 0.15fF
C9 xe inverter_0/A 0.17fF
C10 Nin Oin 0.12fF
C11 Ain bin 0.10fF
C12 VP inverter_0/A 1.64fF
C13 Lin Min 0.12fF
C14 Din Cin 0.10fF
C15 Ein Fin 0.10fF
C16 Pin Oin 0.12fF
C17 Ain VN 0.22fF
C18 bin VN 0.22fF
C19 Cin VN 0.22fF
C20 Din VN 0.22fF
C21 Ein VN 0.22fF
C22 Fin VN 0.22fF
C23 Gin VN 0.22fF
C24 Hin VN 0.22fF
C25 inverter_0/A VN -0.68fF
C26 a_n140_n60# VN -0.14fF
C27 xe VN 1.17fF
C28 inverter_3/a_n10_n20# VN 0.34fF
C29 VP VN 4.95fF
C30 reset_loop VN -1.13fF
C31 inverter_2/A VN 1.62fF
.ends


* Top level circuit neuron

Xpg17Input8p8n_para_1n_0 pg17Input8p8n_para_1n_0/Ain pg17Input8p8n_para_1n_0/bin pg17Input8p8n_para_1n_1/VP
+ pg17Input8p8n_para_1n_0/Din pg17Input8p8n_para_1n_0/Ein pg17Input8p8n_para_1n_0/Fin
+ pg17Input8p8n_para_1n_0/Gin pg17Input8p8n_para_1n_0/Hin pg17Input8p8n_para_1n_0/Cin
+ pg17Input8p8n_para_1n_0/Iin SUB pg17Input8p8n_para_1n_0/Jin pg17Input8p8n_para_1n_0/Kin
+ pg17Input8p8n_para_1n_0/Lin pg17Input8p8n_para_1n_0/Min pg17Input8p8n_para_1n_0/Nin
+ pg17Input8p8n_para_1n_0/Oin pg17Input8p8n_para_1n_0/Pin pg17Input8p8n_para_1n_0/inverter_3/a_n10_n20#
+ pg17Input8p8n_para_1n_0/xe li_n15_275# pg17Input8p8n_para_1n_0/reset_loop pg17Input8p8n_para_1n_0/inverter_2/A
+ pg17Input8p8n_para_1n
Xpg17Input8p8n_para_1n_1 pg17Input8p8n_para_1n_1/Ain pg17Input8p8n_para_1n_1/bin pg17Input8p8n_para_1n_1/VP
+ pg17Input8p8n_para_1n_1/Din pg17Input8p8n_para_1n_1/Ein pg17Input8p8n_para_1n_1/Fin
+ pg17Input8p8n_para_1n_1/Gin pg17Input8p8n_para_1n_1/Hin pg17Input8p8n_para_1n_1/Cin
+ pg17Input8p8n_para_1n_1/Iin SUB pg17Input8p8n_para_1n_1/Jin pg17Input8p8n_para_1n_1/Kin
+ pg17Input8p8n_para_1n_1/Lin pg17Input8p8n_para_1n_1/Min pg17Input8p8n_para_1n_1/Nin
+ pg17Input8p8n_para_1n_1/Oin pg17Input8p8n_para_1n_1/Pin li_n15_275# pg17Input8p8n_para_1n_1/xe
+ pg17Input8p8n_para_1n_1/a_n140_n60# pg17Input8p8n_para_1n_1/reset_loop pg17Input8p8n_para_1n_1/inverter_2/A
+ pg17Input8p8n_para_1n
C0 pg17Input8p8n_para_1n_1/VP li_n15_275# 0.39fF
C1 pg17Input8p8n_para_1n_1/reset_loop pg17Input8p8n_para_1n_0/reset_loop 0.22fF
C2 pg17Input8p8n_para_1n_1/Ain SUB 0.22fF
C3 pg17Input8p8n_para_1n_1/bin SUB 0.22fF
C4 pg17Input8p8n_para_1n_1/Cin SUB 0.22fF
C5 pg17Input8p8n_para_1n_1/Din SUB 0.22fF
C6 pg17Input8p8n_para_1n_1/Ein SUB 0.22fF
C7 pg17Input8p8n_para_1n_1/Fin SUB 0.22fF
C8 pg17Input8p8n_para_1n_1/Gin SUB 0.22fF
C9 pg17Input8p8n_para_1n_1/Hin SUB 0.22fF
C10 pg17Input8p8n_para_1n_1/inverter_0/A SUB -0.82fF
C11 pg17Input8p8n_para_1n_1/a_n140_n60# SUB -0.14fF
C12 pg17Input8p8n_para_1n_1/xe SUB 0.48fF
C13 li_n15_275# SUB 1.92fF
C14 pg17Input8p8n_para_1n_1/reset_loop SUB -1.13fF
C15 pg17Input8p8n_para_1n_1/inverter_2/A SUB 1.53fF
C16 pg17Input8p8n_para_1n_0/Ain SUB 0.22fF
C17 pg17Input8p8n_para_1n_0/bin SUB 0.22fF
C18 pg17Input8p8n_para_1n_0/Cin SUB 0.22fF
C19 pg17Input8p8n_para_1n_0/Din SUB 0.22fF
C20 pg17Input8p8n_para_1n_0/Ein SUB 0.22fF
C21 pg17Input8p8n_para_1n_0/Fin SUB 0.22fF
C22 pg17Input8p8n_para_1n_0/Gin SUB 0.22fF
C23 pg17Input8p8n_para_1n_0/Hin SUB 0.22fF
C24 pg17Input8p8n_para_1n_0/inverter_0/A SUB -0.82fF
C25 pg17Input8p8n_para_1n_0/xe SUB 0.98fF
C26 pg17Input8p8n_para_1n_0/inverter_3/a_n10_n20# SUB 0.34fF
C27 pg17Input8p8n_para_1n_1/VP SUB 8.85fF
C28 pg17Input8p8n_para_1n_0/reset_loop SUB -1.13fF
C29 pg17Input8p8n_para_1n_0/inverter_2/A SUB 1.60fF
.end

