magic
tech sky130A
timestamp 1632866290
<< error_p >>
rect 1048 290 1055 310
rect 1065 273 1072 310
rect 2348 290 2355 310
rect 2365 273 2372 310
rect 3648 290 3655 310
rect 3665 273 3672 310
rect 6248 290 6255 310
rect 6265 273 6272 310
rect 7548 290 7555 310
rect 7565 273 7572 310
rect 8848 290 8855 310
rect 8865 273 8872 310
rect 10148 290 10155 310
rect 10165 273 10172 310
<< error_s >>
rect 4948 290 4955 310
rect 4965 273 4972 310
use 4xpg16in8p8n  4xpg16in8p8n_1 /neural-stationary/Layout
timestamp 1632866290
transform 1 0 5200 0 1 0
box 0 0 5200 755
use 4xpg16in8p8n  4xpg16in8p8n_0
timestamp 1632866290
transform 1 0 0 0 1 0
box 0 0 5200 755
<< end >>
