magic
tech sky130A
timestamp 1632940244
<< poly >>
rect 780 1040 890 1055
rect 875 780 890 1040
rect 875 770 915 780
rect 875 750 885 770
rect 905 750 915 770
rect 875 740 915 750
rect 550 715 590 725
rect 550 695 560 715
rect 580 695 590 715
rect 550 685 590 695
rect 875 520 890 740
rect 860 500 890 520
rect 860 325 875 500
rect 835 315 875 325
rect 755 305 795 315
rect 755 285 765 305
rect 785 285 795 305
rect 835 295 845 315
rect 865 295 875 315
rect 835 285 875 295
rect 755 275 795 285
<< polycont >>
rect 885 750 905 770
rect 560 695 580 715
rect 765 285 785 305
rect 845 295 865 315
<< locali >>
rect -15 1355 880 1375
rect -15 295 5 1355
rect 1051 1200 1066 1220
rect 125 1155 165 1195
rect 190 1155 230 1195
rect 255 1155 295 1195
rect 320 1155 360 1195
rect 385 1155 425 1195
rect 450 1155 490 1195
rect 515 1155 555 1195
rect 580 1155 620 1195
rect 95 785 135 825
rect 160 785 200 825
rect 225 785 265 825
rect 290 785 330 825
rect 355 785 395 825
rect 420 785 460 825
rect 485 785 525 825
rect 550 785 590 825
rect 875 770 915 780
rect 875 750 885 770
rect 905 750 915 770
rect 875 740 915 750
rect 95 685 135 725
rect 160 685 200 725
rect 225 685 265 725
rect 290 685 330 725
rect 355 685 395 725
rect 420 685 460 725
rect 485 685 525 725
rect 550 715 590 725
rect 550 695 560 715
rect 580 695 590 715
rect 550 685 590 695
rect 125 315 165 355
rect 190 315 230 355
rect 255 315 295 355
rect 320 315 360 355
rect 385 315 425 355
rect 450 315 490 355
rect 515 315 555 355
rect 580 315 620 355
rect 1052 350 1096 370
rect 835 315 880 325
rect 755 305 795 315
rect 755 295 765 305
rect -15 285 765 295
rect 785 285 795 305
rect 835 295 845 315
rect 865 310 880 315
rect 865 295 875 310
rect 835 285 875 295
rect 1051 290 1067 310
rect -15 275 795 285
<< metal1 >>
rect 1265 1440 1275 1450
rect 1260 1285 1270 1295
rect 1290 1075 1300 1085
rect 1285 915 1295 925
rect 1285 575 1295 585
rect 1290 425 1300 435
rect 1270 210 1280 220
rect 1265 65 1275 75
use pg17Input8p8n_para_1n  pg17Input8p8n_para_1n_0
timestamp 1632940244
transform 1 0 895 0 1 335
box -930 -335 405 420
use pg17Input8p8n_para_1n  pg17Input8p8n_para_1n_1
timestamp 1632940244
transform 1 0 895 0 -1 1175
box -930 -335 405 420
<< labels >>
rlabel locali -10 750 -10 750 1 ring_loop
rlabel locali 590 325 590 325 1 in1
port 1 n
rlabel locali 525 325 525 325 1 in2
port 2 n
rlabel locali 465 325 465 325 1 in3
port 3 n
rlabel locali 400 330 400 330 1 in4
port 4 n
rlabel locali 330 325 330 325 1 in5
port 5 n
rlabel locali 275 325 275 325 1 in6
port 6 n
rlabel locali 205 335 205 335 1 in7
port 7 n
rlabel locali 145 325 145 325 1 in8
port 8 n
rlabel locali 605 1165 605 1165 1 in9
port 9 n
rlabel locali 520 1160 520 1160 1 in10
port 10 n
rlabel locali 465 1165 465 1165 1 in11
port 11 n
rlabel locali 405 1175 405 1175 1 in12
port 12 n
rlabel locali 335 1160 335 1160 1 in13
port 13 n
rlabel locali 275 1165 275 1165 1 in14
port 14 n
rlabel locali 210 1170 210 1170 1 in15
port 15 n
rlabel locali 145 1170 145 1170 1 in16
port 16 n
rlabel metal1 1270 70 1270 70 1 VP
rlabel metal1 1275 215 1275 215 1 VN
rlabel metal1 1295 430 1295 430 7 VN
rlabel metal1 1290 580 1290 580 1 VP
rlabel locali 510 690 510 690 1 ip2
port 18 n
rlabel locali 435 690 435 690 1 ip3
port 19 n
rlabel locali 380 700 380 700 1 ip4
port 20 n
rlabel locali 305 700 305 700 1 ip5
port 21 n
rlabel locali 240 690 240 690 1 ip6
port 22 n
rlabel locali 180 705 180 705 1 ip7
port 23 n
rlabel locali 105 705 105 705 1 ip8
port 24 n
rlabel locali 565 800 565 800 1 ip9
port 25 n
rlabel locali 500 795 500 795 1 ip10
port 26 n
rlabel locali 435 805 435 805 1 ip11
port 27 n
rlabel locali 370 800 370 800 1 ip12
port 28 n
rlabel locali 305 800 305 800 1 ip13
port 29 n
rlabel locali 240 800 240 800 1 ip14
port 30 n
rlabel locali 175 800 175 800 1 ip15
port 31 n
rlabel locali 110 790 110 790 1 ip16
port 32 n
rlabel metal1 1290 920 1290 920 1 VP
rlabel metal1 1295 1080 1295 1080 7 VN
rlabel metal1 1265 1290 1265 1290 1 VN
port 34 n
rlabel metal1 1270 1445 1270 1445 1 VP
port 33 n
rlabel locali 550 685 590 725 7 Iin
port 14 w
rlabel locali 565 695 565 695 1 ip1
port 17 n
rlabel locali 875 740 915 780 1 ring_loop_branch
port 35 n
<< end >>
