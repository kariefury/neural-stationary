
*PulseLoop
.include sky130nm.lib

Xpg out2 sNoise sNoise sNoise out pg4
Xpg2 out sNoise sNoise sNoise out2 pg4


v2 sNoise  0 dc 0 trrandom (2 20p 0 0.1 .8)
v3 B 0 0.0

.control
tran 0.1ns 10ns
plot v(out2)+4 v(out) v(sNoise)+2
.endc


*PG
.subckt pg4 A B Ap Bp x

xm1 1 reset_loop critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n

xm2 0 A critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm10 0 B critical_node 0 sky130_fd_pr__nfet_01v8 l=150n w=360n
xm11 1 Ap critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm12 1 Bp critical_node 1 sky130_fd_pr__pfet_01v8 l=150n w=720n

xm3 1 critical_node invO 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm4 0 critical_node invO 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm4 1 invO reset_loop 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm5 0 invO reset_loop 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm6 1 invO xe 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm7 0 invO xe 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

xm8 1 xe x 1 sky130_fd_pr__pfet_01v8 l=150n w=720n
xm9 0 xe x 0 sky130_fd_pr__nfet_01v8 l=150n w=360n

v1 1 0 1.8

.ends pg4
