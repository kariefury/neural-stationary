* SPICE3 file created from pg9Input1p8n.ext - technology: sky130A
.include sky130nm.lib
.option scale=10n

Xpg Clk Clk 1 Clk Clk Clk Clk Clk Clk 1 0 out pg9Input1p8n

v2 Clk 0 dc 0 trrandom(2 200p 0 1.9 0.1)
*v2 Clk 0 PULSE 0 1.8 1n 20p 20p 180p 4ns
v1 1 0 1.8

.control
tran 0.1ns 10ns
gnuplot gp v(out) v(Clk)
.endc

.subckt inverter A Y w_n145_115# a_n125_n20#
X0 Y A w_n145_115# w_n145_115# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X1 Y A a_n125_n20# a_n125_n20# sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
.ends

.subckt pg9Input1p8n Ain Bin VP Din Ein Fin Gin Hin Cin Iin VN xout
Xinverter_0 inverter_0/A inverter_2/A VP VN inverter
Xinverter_1 inverter_2/A reset_loop VP VN inverter
Xinverter_2 inverter_2/A xe VP VN inverter
Xinverter_3 xe xout VP VN inverter
X0 a_n390_30# Ein a_n455_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X1 inverter_0/A reset_loop VP VP sky130_fd_pr__pfet_01v8 ad=-0 pd=0 as=0 ps=0 w=100 l=15
X2 a_n585_30# Hin VN VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X3 inverter_0/A Iin VP VP sky130_fd_pr__pfet_01v8 ad=-0 pd=0 as=0 ps=0 w=100 l=15
X4 a_n520_30# Gin a_n585_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X5 a_n195_30# Bin a_n260_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X6 inverter_0/A Ain a_n195_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X7 a_n325_30# Din a_n390_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X8 a_n260_30# Cin a_n325_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X9 a_n455_30# Fin a_n520_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
C0 VP VN 4.21fF
C1 inverter_2/A VN 1.60fF
C2 reset_loop VN -1.07fF
.ends

