* SPICE3 file created from riedelxor2_cyclic.ext - technology: sky130A

X0 xor2_0/a_470_297# xor2_1/B xor2_1/VPWR xor2_0/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X1 xor2_1/VPWR xor2_1/B xor2_0/a_470_297# xor2_0/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 xor2_0/a_112_47# xor2_1/X xor2_1/VGND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X3 xor2_0/a_470_47# xor2_1/X xor2_0/X SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X4 xor2_1/VGND xor2_1/B xor2_0/a_112_47# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X5 xor2_0/a_112_47# xor2_1/B xor2_1/VGND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X6 xor2_1/VGND xor2_1/X xor2_0/a_112_47# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X7 xor2_1/VPWR xor2_1/B xor2_0/a_27_297# xor2_0/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 xor2_0/a_470_297# xor2_1/X xor2_1/VPWR xor2_0/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 xor2_0/X xor2_0/a_112_47# xor2_1/VGND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X10 xor2_1/VPWR xor2_1/X xor2_0/a_470_297# xor2_0/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 xor2_1/VGND xor2_0/a_112_47# xor2_0/X SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X12 xor2_1/VGND xor2_1/B xor2_0/a_470_47# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X13 xor2_0/a_27_297# xor2_1/X xor2_0/a_112_47# xor2_0/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 xor2_0/X xor2_0/a_112_47# xor2_0/a_470_297# xor2_0/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 xor2_0/a_470_297# xor2_0/a_112_47# xor2_0/X xor2_0/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 xor2_0/X xor2_1/X xor2_0/a_470_47# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X17 xor2_0/a_112_47# xor2_1/X xor2_0/a_27_297# xor2_0/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 xor2_0/a_27_297# xor2_1/B xor2_1/VPWR xor2_0/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 xor2_0/a_470_47# xor2_1/B xor2_1/VGND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X20 xor2_1/a_470_297# xor2_1/A xor2_1/VPWR xor2_1/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 xor2_1/VPWR xor2_1/A xor2_1/a_470_297# xor2_1/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X22 xor2_1/a_112_47# xor2_1/B xor2_1/VGND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X23 xor2_1/a_470_47# xor2_1/B xor2_1/X SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X24 xor2_1/VGND xor2_1/A xor2_1/a_112_47# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X25 xor2_1/a_112_47# xor2_1/A xor2_1/VGND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X26 xor2_1/VGND xor2_1/B xor2_1/a_112_47# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X27 xor2_1/VPWR xor2_1/A xor2_1/a_27_297# xor2_1/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 xor2_1/a_470_297# xor2_1/B xor2_1/VPWR xor2_1/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X29 xor2_1/X xor2_1/a_112_47# xor2_1/VGND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X30 xor2_1/VPWR xor2_1/B xor2_1/a_470_297# xor2_1/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 xor2_1/VGND xor2_1/a_112_47# xor2_1/X SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X32 xor2_1/VGND xor2_1/A xor2_1/a_470_47# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X33 xor2_1/a_27_297# xor2_1/B xor2_1/a_112_47# xor2_1/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 xor2_1/X xor2_1/a_112_47# xor2_1/a_470_297# xor2_1/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 xor2_1/a_470_297# xor2_1/a_112_47# xor2_1/X xor2_1/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 xor2_1/X xor2_1/B xor2_1/a_470_47# SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
X37 xor2_1/a_112_47# xor2_1/B xor2_1/a_27_297# xor2_1/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 xor2_1/a_27_297# xor2_1/A xor2_1/VPWR xor2_1/VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 xor2_1/a_470_47# xor2_1/A xor2_1/VGND SUB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=650000u l=150000u
