magic
tech sky130A
magscale 1 2
timestamp 1644013847
<< poly >>
rect 160 681 234 698
rect 160 647 183 681
rect 217 647 234 681
rect 160 616 234 647
rect 3348 643 3432 658
rect 160 518 204 616
rect 3348 609 3375 643
rect 3409 609 3432 643
rect 3348 578 3432 609
rect 3372 264 3410 578
rect 3364 206 3424 264
rect 776 -42 824 24
rect 784 -330 816 -42
rect 2486 -94 2678 -56
rect 756 -347 840 -330
rect 756 -381 783 -347
rect 817 -381 840 -347
rect 756 -412 840 -381
<< polycont >>
rect 183 647 217 681
rect 3375 609 3409 643
rect 783 -381 817 -347
<< locali >>
rect 160 681 234 698
rect 160 647 183 681
rect 217 658 234 681
rect 217 647 3432 658
rect 160 643 3432 647
rect 160 610 3375 643
rect 3346 609 3375 610
rect 3409 609 3432 643
rect 3346 576 3432 609
rect 1162 146 1868 186
rect 1826 132 1868 146
rect 1826 86 2490 132
rect 2448 -96 2490 86
rect 3758 -114 3892 -62
rect 760 -347 834 -330
rect 760 -381 783 -347
rect 817 -381 834 -347
rect 760 -384 834 -381
rect 3844 -384 3892 -114
rect 424 -426 3892 -384
<< metal1 >>
rect 1190 496 2020 592
rect 1946 284 2020 496
rect 1946 188 2630 284
rect 1194 -48 2038 48
rect 1910 -260 2038 -48
rect 1910 -356 2596 -260
use xor2  xor2_1
timestamp 1644004558
transform 1 0 2590 0 1 -308
box -38 -48 1234 592
use xor2  xor2_0
timestamp 1644004558
transform 1 0 0 0 1 0
box -38 -48 1234 592
<< labels >>
rlabel locali 522 634 542 648 1 ainput
port 1 n
rlabel locali 1790 160 1810 174 1 binside
port 2 n
rlabel locali 1760 -410 1780 -396 1 ycyclic
port 3 n
rlabel metal1 1858 534 1878 548 1 powin
port 4 n
rlabel metal1 1818 -14 1838 0 1 gndin
port 5 n
<< end >>
