* SPICE3 file created from neuron.ext - technology: sky130A

.option scale=10000u

.subckt inverter A w_n145_115# a_n10_n20# a_n125_n20#
X0 a_n10_n20# A w_n145_115# w_n145_115# sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X1 a_n10_n20# A a_n125_n20# a_n125_n20# sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
C0 a_n10_n20# w_n145_115# 0.22fF
C1 A a_n125_n20# 0.53fF
C2 a_n10_n20# a_n125_n20# 0.34fF
C3 w_n145_115# a_n125_n20# 0.59fF
.ends

.subckt pg17Input8p8n_para_1n Ain bin VP Din Ein Fin Gin Hin Cin Iin VN Jin Kin Lin
+ Min Nin Oin Pin inverter_3/a_n10_n20# inverter_2/A xe a_n140_n60# reset_loop
Xinverter_0 inverter_0/A VP inverter_2/A VN inverter
Xinverter_1 inverter_2/A VP reset_loop VN inverter
Xinverter_2 inverter_2/A VP xe VN inverter
Xinverter_3 xe VP inverter_3/a_n10_n20# VN inverter
X0 a_n560_30# Ein a_n625_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X1 inverter_0/A reset_loop VP VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=-0 ps=0 w=100 l=15
X2 inverter_0/A a_n140_n60# VN VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X3 inverter_0/A Min inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X4 a_n755_30# Hin VN VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X5 inverter_0/A Kin inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X6 a_n690_30# Gin a_n755_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X7 inverter_0/A Iin inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X8 inverter_0/A Oin inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X9 a_n365_30# bin a_n430_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X10 inverter_0/A Ain a_n365_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X11 inverter_0/A Jin inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X12 a_n495_30# Din a_n560_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X13 inverter_0/A Pin VP VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=-0 ps=0 w=100 l=15
X14 inverter_0/A Nin inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X15 a_n430_30# Cin a_n495_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X16 inverter_0/A Lin inverter_0/A VP sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
X17 a_n625_30# Fin a_n690_30# VN sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=100 l=15
C0 Hin Gin 0.10fF
C1 bin Cin 0.10fF
C2 Din Cin 0.10fF
C3 Din Ein 0.10fF
C4 Ein Fin 0.10fF
C5 Nin Min 0.12fF
C6 Min Lin 0.12fF
C7 inverter_0/A xe 0.17fF
C8 Oin Pin 0.12fF
C9 inverter_0/A VP 1.64fF
C10 Jin Kin 0.12fF
C11 reset_loop VP 0.15fF
C12 Nin Oin 0.12fF
C13 Gin Fin 0.10fF
C14 bin Ain 0.10fF
C15 Jin Iin 0.12fF
C16 Kin Lin 0.12fF
C17 Ain VN 0.22fF
C18 bin VN 0.22fF
C19 Cin VN 0.22fF
C20 Din VN 0.22fF
C21 Ein VN 0.22fF
C22 Fin VN 0.22fF
C23 Gin VN 0.22fF
C24 Hin VN 0.22fF
C25 inverter_0/A VN -0.64fF
C26 a_n140_n60# VN -0.20fF
C27 inverter_3/a_n10_n20# VN 0.34fF
C28 xe VN 1.16fF
C29 inverter_2/A VN 1.63fF
C30 reset_loop VN -1.11fF
C31 VP VN 4.90fF
.ends

.subckt neuron ip1 ring_loop_branch
Xpg17Input8p8n_para_1n_0 pg17Input8p8n_para_1n_0/Ain pg17Input8p8n_para_1n_0/bin pg17Input8p8n_para_1n_1/VP
+ pg17Input8p8n_para_1n_0/Din pg17Input8p8n_para_1n_0/Ein pg17Input8p8n_para_1n_0/Fin
+ pg17Input8p8n_para_1n_0/Gin pg17Input8p8n_para_1n_0/Hin pg17Input8p8n_para_1n_0/Cin
+ ip1 SUB pg17Input8p8n_para_1n_0/Jin pg17Input8p8n_para_1n_0/Kin pg17Input8p8n_para_1n_0/Lin
+ pg17Input8p8n_para_1n_0/Min pg17Input8p8n_para_1n_0/Nin pg17Input8p8n_para_1n_0/Oin
+ pg17Input8p8n_para_1n_0/Pin ring_loop_branch pg17Input8p8n_para_1n_0/inverter_2/A
+ pg17Input8p8n_para_1n_0/xe ring_loop pg17Input8p8n_para_1n_0/reset_loop pg17Input8p8n_para_1n
Xpg17Input8p8n_para_1n_1 pg17Input8p8n_para_1n_1/Ain pg17Input8p8n_para_1n_1/bin pg17Input8p8n_para_1n_1/VP
+ pg17Input8p8n_para_1n_1/Din pg17Input8p8n_para_1n_1/Ein pg17Input8p8n_para_1n_1/Fin
+ pg17Input8p8n_para_1n_1/Gin pg17Input8p8n_para_1n_1/Hin pg17Input8p8n_para_1n_1/Cin
+ pg17Input8p8n_para_1n_1/Iin SUB pg17Input8p8n_para_1n_1/Jin pg17Input8p8n_para_1n_1/Kin
+ pg17Input8p8n_para_1n_1/Lin pg17Input8p8n_para_1n_1/Min pg17Input8p8n_para_1n_1/Nin
+ pg17Input8p8n_para_1n_1/Oin pg17Input8p8n_para_1n_1/Pin ring_loop pg17Input8p8n_para_1n_1/inverter_2/A
+ pg17Input8p8n_para_1n_1/xe ring_loop_branch pg17Input8p8n_para_1n_1/reset_loop pg17Input8p8n_para_1n
C0 ring_loop pg17Input8p8n_para_1n_1/VP 0.43fF
C1 pg17Input8p8n_para_1n_1/reset_loop ring_loop_branch 0.13fF
C2 ring_loop_branch pg17Input8p8n_para_1n_0/reset_loop 0.11fF
C3 pg17Input8p8n_para_1n_1/reset_loop pg17Input8p8n_para_1n_0/reset_loop 0.22fF
C4 pg17Input8p8n_para_1n_1/Ain SUB 0.22fF
C5 pg17Input8p8n_para_1n_1/bin SUB 0.22fF
C6 pg17Input8p8n_para_1n_1/Cin SUB 0.22fF
C7 pg17Input8p8n_para_1n_1/Din SUB 0.22fF
C8 pg17Input8p8n_para_1n_1/Ein SUB 0.22fF
C9 pg17Input8p8n_para_1n_1/Fin SUB 0.22fF
C10 pg17Input8p8n_para_1n_1/Gin SUB 0.22fF
C11 pg17Input8p8n_para_1n_1/Hin SUB 0.22fF
C12 pg17Input8p8n_para_1n_1/inverter_0/A SUB -0.77fF
C13 ring_loop SUB -1.26fF
C14 pg17Input8p8n_para_1n_1/xe SUB 0.46fF
C15 pg17Input8p8n_para_1n_1/inverter_2/A SUB 1.53fF
C16 pg17Input8p8n_para_1n_1/reset_loop SUB -1.11fF
C17 pg17Input8p8n_para_1n_0/Ain SUB 0.22fF
C18 pg17Input8p8n_para_1n_0/bin SUB 0.22fF
C19 pg17Input8p8n_para_1n_0/Cin SUB 0.22fF
C20 pg17Input8p8n_para_1n_0/Din SUB 0.22fF
C21 pg17Input8p8n_para_1n_0/Ein SUB 0.22fF
C22 pg17Input8p8n_para_1n_0/Fin SUB 0.22fF
C23 pg17Input8p8n_para_1n_0/Gin SUB 0.22fF
C24 pg17Input8p8n_para_1n_0/Hin SUB 0.22fF
C25 ip1 SUB -0.38fF
C26 pg17Input8p8n_para_1n_0/inverter_0/A SUB -0.77fF
C27 ring_loop_branch SUB 0.35fF
C28 pg17Input8p8n_para_1n_0/xe SUB 0.97fF
C29 pg17Input8p8n_para_1n_0/inverter_2/A SUB 1.60fF
C30 pg17Input8p8n_para_1n_0/reset_loop SUB -1.11fF
C31 pg17Input8p8n_para_1n_1/VP SUB 8.71fF
.ends

